module launder_clock(input in, output __output);
    assign __output = in;
endmodule


module unlaunder_clock(input in, output __output);
    assign __output = in;
endmodule
